[{"directBlock1":0,"directBlock2":1,"indirectBlock":2,"size":101,"attributes":511},{"directBlock1":5,"directBlock2":6,"indirectBlock":7,"size":188,"attributes":511},{"directBlock1":12,"directBlock2":13,"indirectBlock":14,"size":86,"attributes":511},{"directBlock1":16,"directBlock2":17,"indirectBlock":18,"size":75,"attributes":511},{"directBlock1":20,"directBlock2":21,"indirectBlock":22,"size":68,"attributes":511},{"directBlock1":24,"directBlock2":25,"indirectBlock":26,"size":119,"attributes":511},{"directBlock1":29,"directBlock2":30,"indirectBlock":31,"size":101,"attributes":511},{"directBlock1":34,"directBlock2":-1,"indirectBlock":-1,"size":10,"attributes":511},{"directBlock1":35,"directBlock2":36,"indirectBlock":37,"size":166,"attributes":511},{"directBlock1":42,"directBlock2":-1,"indirectBlock":-1,"size":1,"attributes":511},null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null,null]