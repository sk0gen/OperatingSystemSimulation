{"blockSize":32,"size":2048,"disk":["M","O","V"," ","A"," ","0",";","\n","M","O","V"," ","B"," ","1",";","\n","M","O","V"," ","C"," ","1","4",";","\n","M","O","V"," ","D"," ","B",";","\n","A","D","D"," ","B"," ","A",";","\n","M","O","V"," ","A"," ","D",";","\n","D","E","C"," ","C",";","\n","J","N","\u0003","\u0004","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","Z"," ","2","5",";","\n","H","L","W"," ","K","o","n","i","e","c",";","\n","P","R","I","N","T","F","L","A","G","S",";","\r","\n","R","E","T"," ","0",";","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","H","L","W"," ","S","t","a","r","t","P","i","p","e","s","1",";","\n","C","P"," ","t","e","s","t","P","i","p","e","s","2",".","a","s","m",";","\n","C","O","P"," ","p","i","p","1"," ","0",";","\n","S","M","P"," ","p","i","p","1"," ","1",";","\n","S","M","P"," ","\b","\t","\n","\u000b","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","p","i","p","1"," ","2",";","\n","S","M","P"," ","p","i","p","1"," ","3",";","\n","S","M","P"," ","p","i","p","1"," ","4",";","\n","S","M","P"," ","p","i","p","1"," ","5",";","\n","S","M","P"," ","p","i","p","1"," ","6",";","\n","S","M","P"," ","p","i","p","1"," ","7",";","\n","S","M","P"," ","p","i","p","1"," ","8",";","\n","S","M","P"," ","p","i","p","1"," ","9",";","\n","D","O","P"," ","p","i","p","1",";","\n","H","L","W"," ","E","n","d","P","i","p","e","s","1",";","\n","R","E","T"," ","0",";","\n","ÿ","ÿ","ÿ","ÿ","H","L","W"," ","S","t","a","r","t","P","i","p","e","s","2",";","\n","M","O","V"," ","B"," ","9",";","\n","R","M","P"," ","p","i","p","1",";","\n","P","O","P"," ","A",";","\n","P","R","T"," ","A",";","\n","D","E","C"," ","B",";","\n","J","N","Z"," ","2","4",";","\u000f","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","\n","H","L","W"," ","E","n","d","P","i","p","e","s","2",";","\n","R","E","T"," ","0",";","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","H","L","W"," ","C","z","e","k","a","m","N","a","W","a","r","u","n","e","k","1",";","\r","\n","C","P"," ","t","e","s","t","C","o","n","d","2",".","a","s","m",";","\r","\n","W","A","T"," ","1",";","\r","\n","H","L","W"," ","P","r","z","e","s","z","e","d","l","e","\u0013","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","m","1",";","\r","\n","R","E","T"," ","0",";","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","H","L","W"," ","S","t","a","r","t","2",";","\n","M","O","V"," ","A"," ","5","0",";","\n","D","E","C"," ","A",";","\n","J","N","Z"," ","2","0",";","\n","H","L","W"," ","i","d","z","i","e","S","y","g","n","a","l","2",";","\n","S","I","G"," ","1",";","\n","R","E","\u0017","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","T"," ","0",";","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","H","L","W"," ","w","c","h","o","d","z","e","D","o","Z","a","m","k","a","1",";","\n","C","P"," ","t","e","s","t","L","o","c","k","2",".","a","s","m",";","\n","M","O","V"," ","A"," ","5","0",";","\n","L","C","K"," ","1",";","\n","D","E","C"," ","A",";","\n","H","\u001b","\u001c","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","L","W"," ","s","i","e","d","z","e","W","Z","a","m","k","u","1",";","\n","J","N","Z"," ","5","2",";","\n","U","N","L"," ","1",";","\n","H","L","W"," ","w","y","s","z","e","d","l","e","m","1",";","\n","R","E","T"," ","0",";","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","H","L","W"," ","w","c","h","o","d","z","e","D","o","Z","a","m","k","a","2",";","\n","M","O","V"," ","A"," ","5","0",";","\n","L","C","K"," ","1",";","\n","D","E","C"," ","A",";","\n","H","L","W"," ","s","i","e","d","z","e","W","Z","a","m","k","u","2",";","\n"," ","!","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","J","N","Z"," ","3","5",";","\n","U","N","L"," ","1",";","\n","H","L","W"," ","w","y","s","z","e","d","l","e","m","2",";","\n","R","E","T"," ","0",";","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","1","2","3","4","5","6","7","8","8","\n","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","H","L","W"," ","o","d","c","z","y","t","_","p","l","i","k","u","_","d","a","n","e",".","t","x","t",";","\n","R","D","F"," ","d","a","n","e",".","t","x","t",";","\n","P","O","P"," ","D",";","\n","P","O","P"," ","A",";","\n","S","U","B"," ","D"," ","1",";","\n","\u0026","\u0027","(",")","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","P","O","P"," ","B",";","\n","A","D","D"," ","A"," ","B",";","\n","D","E","C"," ","D",";","\n","J","N","Z"," ","5","9",";","\n","H","L","W"," ","s","u","m","a",":",";","\n","P","R","T"," ","A",";","\n","R","M","F"," ","w","y","n","i","k",".","t","x","t",";","\n","C","R","F"," ","w","y","n","i","k",".","t","x","t",";","\n","W","R","F"," ","w","y","n","i","k",".","t","x","t"," ","A",";","\n","R","E","T"," ","0",";","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","$","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ","ÿ"]}