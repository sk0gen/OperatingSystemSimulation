{"testPipes2.asm":2,"testPipes1.asm":1,"fib.asm":0,"testCond2.asm":4,"wynik.txt":9,"testLock2.asm":6,"testCond1.asm":3,"testLock1.asm":5,"testDisk.asm":8,"dane.txt":7}